
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY LATCH16 IS
   PORT ( CLK : IN STD_LOGIC;
          I: IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
   		);
END LATCH16;


ARCHITECTURE BEHAVIOR OF LATCH16 IS
SIGNAL SIG: STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
BEGIN     
    O <= SIG;
    	
	WRITE: PROCESS (CLK)
	BEGIN
		IF RISING_EDGE (CLK) THEN
			SIG <= I;	
		END IF;
	END PROCESS WRITE;
	  
END BEHAVIOR;

