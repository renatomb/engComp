
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY CPU_OP IS
	PORT (	CLK_1, CLK_2, CLK_3: 	 		 IN  STD_LOGIC;	-- CLOCKS
			N, Z,											-- SINAIS DE TESTE VINDOS DA ULA
	        OUT_RD, OUT_WR:   				 OUT STD_LOGIC;	-- SINAIS DE CONTROLE P/ MEMORIA
			AMUX, 											-- CONTROLA A ENTRADA ESQUERDA DA ULA
			MBR, 											-- CARREGA MBR A PARTIR DO DESLOCADOR
			MAR, 											-- CARREGA MAR A PARTIR DO LATCH B
			IN_RD, 										    -- REQUISITA LEITURA DA MEM�RIA
			IN_WR,  										-- REQUISITA ESCRITA NA MEM�RIA
			ENC:			  				  IN STD_LOGIC;	-- HABILITA BARRAMENTO C
			ULA, 											-- CONTROLA OPERA��ES DA ULA
			SH:			IN 	STD_LOGIC_VECTOR ( 1 DOWNTO 0);	-- CONTROLA O DESLOCDOR NA SAIDA DA ULA
			A, B,											-- DEFINE ENDERECOS DE LEITURA DOS REGS DA MEM�RIA DE RASCUNHO
			C: 			IN  STD_LOGIC_VECTOR ( 3 DOWNTO 0); -- DEFINE ENDERECOS DE ESCRITA DOS REGS DA MEM�RIA DE RASCUNHO
			ADD_MEM:	OUT STD_LOGIC_VECTOR (11 DOWNTO 0);	-- LIGACAO COM BARRAMENTO DE ENDERECOS 
	        OUT_MEM:	OUT STD_LOGIC_VECTOR (15 DOWNTO 0);	-- LIGACAO COM BARRAMENTO DE DADOS
	         IN_MEM:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0));-- LIGACAO COM BARRAMENTO DE DADOS

END CPU_OP;


ARCHITECTURE BEHAVIOR OF CPU_OP IS

COMPONENT DECOD4_TO_16 IS
   PORT ( I: IN   STD_LOGIC_VECTOR ( 3 DOWNTO 0 );
          O: OUT  STD_LOGIC_VECTOR (15 DOWNTO 0 )
        );
END COMPONENT;

COMPONENT DESLOCADOR16 IS
   PORT ( S: IN  STD_LOGIC_VECTOR ( 1 DOWNTO 0);
          I: IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
END COMPONENT;

COMPONENT MEM_RASCUNHO16x16 IS
   PORT ( CLK: IN STD_LOGIC; 
   		  SA, SB, SC: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
          BAR_C: IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  BAR_A: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  BAR_B: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
END COMPONENT;

COMPONENT LATCH16 IS
   PORT ( CLK: IN STD_LOGIC;
          I: IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
   		);
END COMPONENT;

COMPONENT MUX16_2_TO_1 IS
   PORT ( S:  IN   STD_LOGIC;
   		  I0: IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
          I1: IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
          O:  OUT  STD_LOGIC_VECTOR ( 15 DOWNTO 0 )
        );
END COMPONENT;

COMPONENT REGISTRADOR_D16 IS
   PORT ( CLK, RD_MEM, WR_MEM, RD_CPU: IN STD_LOGIC;
          I_CPU:  IN    STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O_CPU:  OUT   STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  I_MEM:  IN    STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O_MEM:  OUT   STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
END COMPONENT;

COMPONENT REGISTRADOR_E12 IS
   PORT ( CLK, E: IN STD_LOGIC;
          I: IN  STD_LOGIC_VECTOR (11 DOWNTO 0);
   		  O: OUT STD_LOGIC_VECTOR (11 DOWNTO 0)
        );
END COMPONENT;

COMPONENT ULA16 IS
   PORT ( S:   IN   STD_LOGIC_VECTOR (  1 DOWNTO 0 );
          A:   IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
          B:   IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
		  O:   OUT  STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
          N,Z: OUT  STD_LOGIC
        );
END COMPONENT;

SIGNAL BAR_A, BAR_B, BAR_C, SIG_LATCH_A, SIG_LATCH_B,
       SIG_LEFT_ULA, SIG_SHIFT, SIG_LEFT_AMUX,
       SIG_RAS_A, SIG_RAS_B, SIG_RAS_C, SIGT_RAS_C: STD_LOGIC_VECTOR ( 15 DOWNTO 0); 

BEGIN

OUT_RD <= IN_RD;
OUT_WR <= IN_WR;

UNIT_ULA: 
	ULA16
	PORT MAP (ULA, SIG_LEFT_ULA, SIG_LATCH_B, SIG_SHIFT, N, Z);

UNIT_SHIFT:
	DESLOCADOR16
	PORT MAP (SH, SIG_SHIFT, BAR_C);

UNIT_MBR:
	REGISTRADOR_D16
	PORT MAP (CLK_3, IN_RD, IN_WR, MBR, BAR_C, SIG_LEFT_AMUX, IN_MEM, OUT_MEM);

UNIT_MAR:
	REGISTRADOR_E12
	PORT MAP (CLK_2, MAR, SIG_LATCH_B(11 DOWNTO 0), ADD_MEM);

UNIT_AMUX:
	MUX16_2_TO_1
	PORT MAP (AMUX, SIG_LATCH_A, SIG_LEFT_AMUX, SIG_LEFT_ULA);

UNIT_LATCH_A:
	LATCH16
	PORT MAP (CLK_1, BAR_A, SIG_LATCH_A);

UNIT_LATCH_B:
	LATCH16
	PORT MAP (CLK_1, BAR_B, SIG_LATCH_B);

UNIT_REGS:
	MEM_RASCUNHO16x16
	PORT MAP (CLK_3, SIG_RAS_A, SIG_RAS_B, SIG_RAS_C, BAR_C, BAR_A, BAR_B);

UNIT_DECOD_A:
	DECOD4_TO_16 
	PORT MAP (A, SIG_RAS_A);

UNIT_DECOD_B:
	DECOD4_TO_16
	PORT MAP (B, SIG_RAS_B);

UNIT_DECOD_C:
	DECOD4_TO_16
	PORT MAP (C, SIGT_RAS_C);

ENC_END_C:
	FOR I IN 0 TO 15 GENERATE
		SIG_RAS_C(I) <= ENC AND SIGT_RAS_C(I);
	END GENERATE;

END BEHAVIOR;

