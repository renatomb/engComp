

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY ULA16 IS
	PORT ( S:    IN   STD_LOGIC_VECTOR (  1 DOWNTO 0 );     --SELECIONA OPERACAO
           A:    IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );		--OPERANDO A
           B:    IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );		--OPERANDO B
		   O:    OUT  STD_LOGIC_VECTOR ( 15 DOWNTO 0 );	    --RESULTADO
           N,												--RESULTADO DA OPERACAO EH NEGATIVO
           Z: OUT  STD_LOGIC );								--RESULTADO DA OPERACAO EH ZERO
END ULA16;


ARCHITECTURE BEHAVIOR OF ULA16 IS

   SIGNAL SIG_S: STD_LOGIC_VECTOR ( 3 DOWNTO 0 );
   SIGNAL SIG_O: STD_LOGIC_VECTOR (15 DOWNTO 0 );
   SIGNAL SUM:	 STD_LOGIC_VECTOR (15 DOWNTO 0 ); 	

BEGIN

   SIG_S(0) <= (NOT S(0)) AND (NOT S(1));
   SIG_S(1) <= S(0) AND (NOT S(1));
   SIG_S(2) <= (NOT S(0)) AND S(1);
   SIG_S(3) <= S(0) AND S(1);
   
   SUM <= A+B;
  
GEN_SIGNAL_OUT:
	FOR I IN 0 TO 15 GENERATE
		SIG_O(I) <= ((SIG_S(0) AND SUM(I)) OR
					 (SIG_S(1) AND A(I) AND B(I)) OR
                  	 (SIG_S(2) AND A(I)) OR
                  	 (SIG_S(3) AND NOT A(I))); 
	END GENERATE GEN_SIGNAL_OUT;	

OUTPUTS:   
   O <= SIG_O;
   N <= SIG_O(15);
   Z <= NOT (SIG_O(0) OR SIG_O(1) OR SIG_O(2)  OR SIG_O(3)  OR SIG_O(4)  OR SIG_O(5)  OR SIG_O(6)  OR SIG_O(7) OR
        	 SIG_O(8) OR SIG_O(9) OR SIG_O(10) OR SIG_O(11) OR SIG_O(12) OR SIG_O(13) OR SIG_O(14) OR SIG_O(15));
	 
END BEHAVIOR;
