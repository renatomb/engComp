
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY REGISTRADOR_D16 IS
   PORT ( CLK, RD_MEM, WR_MEM, RD_CPU: IN STD_LOGIC;
          I_CPU:  IN    STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O_CPU:  OUT   STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  I_MEM:  IN    STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O_MEM:  OUT   STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
END REGISTRADOR_D16;


ARCHITECTURE BEHAVIOR OF REGISTRADOR_D16 IS
SIGNAL SIG: STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
BEGIN     
    O_CPU <= SIG;
    	
	REG_CHANGE: PROCESS (CLK, RD_MEM, WR_MEM, RD_CPU)
	BEGIN
		IF RISING_EDGE (CLK) THEN
			IF RD_MEM='1' THEN
				SIG <= I_MEM;
			ELSE
				IF RD_CPU='1' THEN
					SIG <= I_CPU;
				END IF;	
				IF WR_MEM='1' THEN
					O_MEM <= I_CPU;
				END IF;
			END IF;				
		END IF;
	END PROCESS REG_CHANGE;
	  
END BEHAVIOR;
