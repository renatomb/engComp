
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY CPU IS
	PORT ( -------------------
	       CLK: IN STD_LOGIC;
	       -------------------	
		   RD, WR:   OUT STD_LOGIC;							-- SINAIS DE CONTROLE P/ MEMORIA
	       ADD_MEM:  OUT STD_LOGIC_VECTOR(11 DOWNTO 0);		-- LIGACAO COM BARRAMENTO DE ENDERECOS 
	       OUT_MEM:  OUT STD_LOGIC_VECTOR(15 DOWNTO 0);		-- DEFINE DADOS DA MEM�RIA
			IN_MEM:  IN  STD_LOGIC_VECTOR(15 DOWNTO 0));	-- DEFINE DADOS DA MEM�RIA
END CPU;


ARCHITECTURE BEHAVIOR OF CPU IS

COMPONENT CPU_CONTROLLER IS
	PORT (	CLK, N, Z: IN STD_LOGIC;
	    	AMUX, MBR,	MAR, RD, WR, ENC: OUT STD_LOGIC;	 							
			ULA, SH:  OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			A, B, C:  OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT CPU_OP IS
	PORT (	CLK_1, CLK_2, CLK_3: IN  STD_LOGIC;	
			N, Z, OUT_RD, OUT_WR: OUT STD_LOGIC;	
			AMUX, MBR, MAR, IN_RD, IN_WR, ENC: IN STD_LOGIC;	
			ULA, SH:		IN 	STD_LOGIC_VECTOR ( 1 DOWNTO 0);	
			A, B, C: 		IN  STD_LOGIC_VECTOR ( 3 DOWNTO 0);  
			ADD_MEM:		OUT STD_LOGIC_VECTOR (11 DOWNTO 0);	
	        OUT_MEM:		OUT STD_LOGIC_VECTOR (15 DOWNTO 0);	
	         IN_MEM:		IN  STD_LOGIC_VECTOR (15 DOWNTO 0));
END COMPONENT;

COMPONENT CLOCK IS
	PORT (	O: OUT STD_LOGIC);
END COMPONENT;

SIGNAL SIG_CLK_1, SIG_CLK_2, SIG_CLK_3, SIG_CLK_4,
       SIG_N, SIG_Z, SIG_AMUX, SIG_MBR, SIG_MAR, SIG_RD, SIG_WR, SIG_ENC : STD_LOGIC;
SIGNAL SIG_ULA, SIG_SH: STD_LOGIC_VECTOR(1 DOWNTO 0); 			
SIGNAL SIG_A, SIG_B, SIG_C: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL SIG_COUNT: STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN

CONTROLLER:
    CPU_CONTROLLER
    PORT MAP (SIG_CLK_1, SIG_N, SIG_Z,
    		  SIG_AMUX, SIG_MBR, SIG_MAR, SIG_RD, SIG_WR, SIG_ENC, 
    		  SIG_ULA, SIG_SH,
    		  SIG_A, SIG_B, SIG_C);
OPERATOR:    						 
    CPU_OP
    PORT MAP (SIG_CLK_2, SIG_CLK_3, SIG_CLK_4,
              SIG_N, SIG_Z, RD, WR,
              SIG_AMUX, SIG_MBR, SIG_MAR, SIG_RD, SIG_WR, SIG_ENC, 
      		  SIG_ULA, SIG_SH,
    		  SIG_A, SIG_B, SIG_C,
    		  ADD_MEM,
              OUT_MEM,
              IN_MEM);

COUNTER:
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE (CLK) THEN
			CASE SIG_COUNT IS
				WHEN "00" => SIG_COUNT <= "01";
				WHEN "01" => SIG_COUNT <= "10";
				WHEN "10" => SIG_COUNT <= "11";
				WHEN "11" => SIG_COUNT <= "00";
				WHEN OTHERS =>
			END CASE;
		END IF;
	END PROCESS COUNTER;
			
GEN_CLKS:
	PROCESS (SIG_COUNT)
	BEGIN
		IF SIG_COUNT = "00" THEN
			SIG_CLK_1 <= '1';
			--SIG_CLK_2 <= '0';
	        --SIG_CLK_3 <= '0';
	        SIG_CLK_4 <= '0';
		ELSIF SIG_COUNT = "01" THEN
			SIG_CLK_1 <= '0';
			SIG_CLK_2 <= '1';
	        --SIG_CLK_3 <= '0';
	        --SIG_CLK_4 <= '0';	
		ELSIF SIG_COUNT = "10" THEN
			--SIG_CLK_1 <= '0';
			SIG_CLK_2 <= '0';
	        SIG_CLK_3 <= '1';
	        --SIG_CLK_4 <= '0';
		ELSE
			--SIG_CLK_1 <= '0';
			--SIG_CLK_2 <= '0';
	        SIG_CLK_3 <= '0';
	        SIG_CLK_4 <= '1';
		END IF;
	END PROCESS GEN_CLKS;					 	
				
END BEHAVIOR;

