
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY MEM_RASCUNHO16x16 IS
   PORT ( CLK: IN STD_LOGIC; 
   		  SA, SB, SC: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
          BAR_C: IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
   		  BAR_A: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
   		  BAR_B: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
        );
END MEM_RASCUNHO16x16;


ARCHITECTURE BEHAVIOR OF MEM_RASCUNHO16x16 IS

SUBTYPE REG IS STD_LOGIC_VECTOR( 15 DOWNTO 0 );
TYPE REGS IS ARRAY (15 DOWNTO 0) OF REG;
SIGNAL SIG: REGS;

BEGIN

	SIG(5)<="0000000000000000";
	SIG(6)<="0000000000000001";
	SIG(7)<="1000000000000001";
	SIG(8)<="0000111111111111";
	SIG(9)<="0000000011111111";
	      
	REG_WRITE_C: PROCESS (CLK, SC)
	BEGIN
		IF RISING_EDGE (CLK) THEN
			CASE SC IS
				WHEN "0000000000000001" => SIG(0) <= BAR_C;
				WHEN "0000000000000010" => SIG(1) <= BAR_C;
				WHEN "0000000000000100" => SIG(2) <= BAR_C;
				WHEN "0000000000001000" => SIG(3) <= BAR_C;
				WHEN "0000000000010000" => SIG(4) <= BAR_C;
				WHEN "0000010000000000" => SIG(10) <= BAR_C;
				WHEN "0000100000000000" => SIG(11) <= BAR_C;
				WHEN "0001000000000000" => SIG(12) <= BAR_C;
				WHEN "0010000000000000" => SIG(13) <= BAR_C;
				WHEN "0100000000000000" => SIG(14) <= BAR_C;
				WHEN "1000000000000000" => SIG(15) <= BAR_C;
				WHEN OTHERS =>
			END CASE;
		END IF;
	END PROCESS REG_WRITE_C;
	
    REG_READ_A: PROCESS (SA)
	BEGIN
		--IF RISING_EDGE (CLK) THEN
			CASE SA IS
				WHEN "0000000000000001" => BAR_A <= SIG(0);
				WHEN "0000000000000010" => BAR_A <= SIG(1);
				WHEN "0000000000000100" => BAR_A <= SIG(2);
				WHEN "0000000000001000" => BAR_A <= SIG(3);
				WHEN "0000000000010000" => BAR_A <= SIG(4);
				WHEN "0000000000100000" => BAR_A <= SIG(5);
				WHEN "0000000001000000" => BAR_A <= SIG(6);
				WHEN "0000000010000000" => BAR_A <= SIG(7);
				WHEN "0000000100000000" => BAR_A <= SIG(8);
				WHEN "0000001000000000" => BAR_A <= SIG(9);
				WHEN "0000010000000000" => BAR_A <= SIG(10);
				WHEN "0000100000000000" => BAR_A <= SIG(11);
				WHEN "0001000000000000" => BAR_A <= SIG(12);
				WHEN "0010000000000000" => BAR_A <= SIG(13);
				WHEN "0100000000000000" => BAR_A <= SIG(14);
				WHEN "1000000000000000" => BAR_A <= SIG(15);
				WHEN OTHERS =>
			END CASE;
		--END IF;
	END PROCESS REG_READ_A;
	
	REG_READ_B: PROCESS (SB)
	BEGIN
		--IF RISING_EDGE (CLK) THEN
			CASE SB IS
				WHEN "0000000000000001" => BAR_B <= SIG(0);
				WHEN "0000000000000010" => BAR_B <= SIG(1);
				WHEN "0000000000000100" => BAR_B <= SIG(2);
				WHEN "0000000000001000" => BAR_B <= SIG(3);
				WHEN "0000000000010000" => BAR_B <= SIG(4);
				WHEN "0000000000100000" => BAR_B <= SIG(5);
				WHEN "0000000001000000" => BAR_B <= SIG(6);
				WHEN "0000000010000000" => BAR_B <= SIG(7);
				WHEN "0000000100000000" => BAR_B <= SIG(8);
				WHEN "0000001000000000" => BAR_B <= SIG(9);
				WHEN "0000010000000000" => BAR_B <= SIG(10);
				WHEN "0000100000000000" => BAR_B <= SIG(11);
				WHEN "0001000000000000" => BAR_B <= SIG(12);
				WHEN "0010000000000000" => BAR_B <= SIG(13);
				WHEN "0100000000000000" => BAR_B <= SIG(14);
				WHEN "1000000000000000" => BAR_B <= SIG(15);
				WHEN OTHERS =>
			END CASE;
		--END IF;
	END PROCESS REG_READ_B;
	  
END BEHAVIOR;

