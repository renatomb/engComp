

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY DESLOCADOR16 IS
   PORT ( S: IN  STD_LOGIC_VECTOR ( 1 DOWNTO 0);
          I: IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
   		  O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
END DESLOCADOR16;


ARCHITECTURE BEHAVIOR OF DESLOCADOR16 IS
BEGIN
  
	DO_SHIFT: PROCESS (I,S)
	BEGIN
		CASE S IS
				WHEN "01" => O <= I(14 DOWNTO 0) & '0';
				WHEN "10" => O <= '0' & I(15 DOWNTO 1) ;
				WHEN OTHERS => O <= I;	
    	END CASE;		
	END PROCESS DO_SHIFT;
	  
END BEHAVIOR;
