
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY REGISTRADOR_E12 IS
   PORT ( CLK, E: IN STD_LOGIC;
          I: IN  STD_LOGIC_VECTOR (11 DOWNTO 0);
   		  O: OUT STD_LOGIC_VECTOR (11 DOWNTO 0)
   		);
END REGISTRADOR_E12;


ARCHITECTURE BEHAVIOR OF REGISTRADOR_E12 IS
SIGNAL SIG: STD_LOGIC_VECTOR ( 11 DOWNTO 0 );
BEGIN     
    O <= SIG;
    	
	REG_WRITE: PROCESS (CLK, E)
	BEGIN
		IF RISING_EDGE (CLK) THEN
			IF E='1' THEN
				SIG <= I;	
			END IF;		
		END IF;
	END PROCESS REG_WRITE;
	  
END BEHAVIOR;
