
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY MUX16_2_TO_1 IS
   PORT ( S:  IN   STD_LOGIC;
   		  I0: IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
          I1: IN   STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
          O:  OUT  STD_LOGIC_VECTOR ( 15 DOWNTO 0 ));
END MUX16_2_TO_1;


ARCHITECTURE BEHAVIOR OF MUX16_2_TO_1 IS
BEGIN
   WITH S SELECT
     O <= I0 WHEN '0',
          I1 WHEN OTHERS;  
END BEHAVIOR;
